LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Timer IS
PORT (
	Clk : IN STD_LOGIC;
	Sel_Switch : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
	Reset_N : IN STD_LOGIC;
	Hex2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	Hex1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	Hex0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
	Test : OUT STD_LOGIC
);
END Timer;

ARCHITECTURE arch OF Timer IS

BEGIN

